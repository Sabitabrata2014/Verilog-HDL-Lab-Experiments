module or_m (p,q,r);

input p,q;
output r;

assign r=p | q;

endmodule