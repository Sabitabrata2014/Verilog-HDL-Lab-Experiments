`timescale 1ns / 1ps

module tff_m_tb; 

reg t; 
reg rst;
reg clk;

wire q;
wire qbar; 

tff_m DUT(t,rst,clk,q,qbar); 

always begin
#20 clk=~clk;
end

initial begin 

clk=1'b0;
t=1'b0;
rst=1'b1;#100;

rst=1'b0;

t=1'b1;#80;
t=1'b0;#120;
t=1'b1;#100;

end 
endmodule 